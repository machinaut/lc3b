// alu.vh - ALU header file

`ifndef _alu_vh_
`define _alu_vh_

// ALU operations
`define ALUK_ADD   2'b00 // A + B
`define ALUK_AND   2'b01 // A & B
`define ALUK_XOR   2'b10 // A ^ B
`define ALUK_PASSA 2'b11 // A

`endif //_alu_vh_
